**************24CLK_divider_CMOS*************
.subckt clkdivider N001 0 N008 Q4
XU1 0 N001 N003 0 0 Q0 N003 N008 DFFSR
XU2 0 N001 N004 0 0 Q1 N004 N003 DFFSR
XU3 0 N001 N005 0 0 Q2 N005 N004 DFFSR
XU4 0 N001 N006 0 N002 Q3 N006 Q2 DFFSR
XU5 0 N001 N007 0 N002 Q4 N007 N006 DFFSR
XU6 N001 0 Q3 Q4 N002 AND
.ends clkdivider

**********DFF*************
.subckt DFFSR 0 1 D S_ R_ Q Q_bar CLK
Msp S S_ 1 1 pfet w=2u l=0.2u
Msn S S_ 0 0 nfet w=1u l=0.2u
Mrp R R_ 1 1 pfet w=2u l=0.2u
Mrn R R_ 0 0 nfet w=1u l=0.2u
M0 a R 1 1 pfet w=2u l=0.2u
M1 1 b a 1 pfet w=2u l=0.2u
M2 b c 1 1 pfet w=2u l=0.2u
M3 1 S b 1 pfet w=2u l=0.2u
M4 c dd a 1 pfet w=1u l=0.2u
M5 e f c 1 pfet w=1u l=0.2u
M6 1 D e 1 pfet w=2u l=0.2u
M7 1 dd f 1 pfet w=2u l=0.2u
M8 dd CLK 1 1 pfet w=2u l=0.2u
M9 g dd b 1 pfet w=1u l=0.2u
M10 h f g 1 pfet w=1u l=0.2u
M11 Q_bar g 1 1 pfet w=2u l=0.2u
M12 1 R Q_bar 1 pfet w=2u l=0.2u
M13 h Q_bar 1 1 pfet w=2u l=0.2u
M14 1 S h 1 pfet w=2u l=0.2u
M15 1 Q_bar Q 1 pfet w=2u l=0.2u
M16 j R a 0 nfet w=2u l=0.2u
M17 0 b j 0 nfet w=2u l=0.2u
M18 k c 0 0 nfet w=2u l=0.2u
M19 b S k 0 nfet w=2u l=0.2u
M20 c f a 0 nfet w=1u l=0.2u
M21 e dd c 0 nfet w=1u l=0.2u
M22 0 D e 0 nfet w=1u l=0.2u
M23 0 dd f 0 nfet w=1u l=0.2u
M24 dd CLK 0 0 nfet w=1u l=0.2u
M25 g f b 0 nfet w=1u l=0.2u
M26 h dd g 0 nfet w=1u l=0.2u
M27 l g Q_bar 0 nfet w=2u l=0.2u
M28 0 R l 0 nfet w=2u l=0.2u
M29 m Q_bar 0 0 nfet w=2u l=0.2u
M30 h S m 0 nfet w=2u l=0.2u
M31 0 Q_bar Q 0 nfet w=1u l=0.2u
.ends DFFSR

*****AND*****

.subckt AND N001 0 N003 N004 OUT
M1 N001 N003 N002 N001 pfet l=0.2u w=2u
M2 N001 N004 N002 N001 pfet l=0.2u w=2u
M3 N002 N003 N005 0 nfet l=0.2u w=1u
M5 N001 N002 OUT N001 pfet l=0.2u w=2u
M6 OUT N002 0 0 nfet l=0.2u w=1u
M4 N005 N004 0 0 nfet l=0.2u w=1u
.ends AND


X1 1_d 0 clk clk1 clkdivider 

************************************
.include osu018.lib

************************************

Vdda 1_d 0 1.8
Vclk clk 0 pulse(0 1.8 1n 1n 1n 0.25u 0.5u)


.tran 1u 30u
.control
run
plot V(clk1) V(clk)
.endc
.end
