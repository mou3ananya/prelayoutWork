******CLK_DIVIDER*************

.inc osu018.lib


*******************DFFSR***********************

.subckt DFFSR 0 1 D S_ R_ Q Q_bar CLK
Msp S S_ 1 1 pfet w=2u l=0.2u
Msn S S_ 0 0 nfet w=1u l=0.2u
Mrp R R_ 1 1 pfet w=2u l=0.2u
Mrn R R_ 0 0 nfet w=1u l=0.2u
M0 a R 1 1 pfet w=2u l=0.2u
M1 1 b a 1 pfet w=2u l=0.2u
M2 b c 1 1 pfet w=2u l=0.2u
M3 1 S b 1 pfet w=2u l=0.2u
M4 c dd a 1 pfet w=1u l=0.2u
M5 e f c 1 pfet w=1u l=0.2u
M6 1 D e 1 pfet w=2u l=0.2u
M7 1 dd f 1 pfet w=2u l=0.2u
M8 dd CLK 1 1 pfet w=2u l=0.2u
M9 g dd b 1 pfet w=1u l=0.2u
M10 h f g 1 pfet w=1u l=0.2u
M11 Q_bar g 1 1 pfet w=2u l=0.2u
M12 1 R Q_bar 1 pfet w=2u l=0.2u
M13 h Q_bar 1 1 pfet w=2u l=0.2u
M14 1 S h 1 pfet w=2u l=0.2u
M15 1 Q_bar Q 1 pfet w=2u l=0.2u
M16 j R a 0 nfet w=2u l=0.2u
M17 0 b j 0 nfet w=2u l=0.2u
M18 k c 0 0 nfet w=2u l=0.2u
M19 b S k 0 nfet w=2u l=0.2u
M20 c f a 0 nfet w=1u l=0.2u
M21 e dd c 0 nfet w=1u l=0.2u
M22 0 D e 0 nfet w=1u l=0.2u
M23 0 dd f 0 nfet w=1u l=0.2u
M24 dd CLK 0 0 nfet w=1u l=0.2u
M25 g f b 0 nfet w=1u l=0.2u
M26 h dd g 0 nfet w=1u l=0.2u
M27 l g Q_bar 0 nfet w=2u l=0.2u
M28 0 R l 0 nfet w=2u l=0.2u
M29 m Q_bar 0 0 nfet w=2u l=0.2u
M30 h S m 0 nfet w=2u l=0.2u
M31 0 Q_bar Q 0 nfet w=1u l=0.2u
.ends DFFSR


****************AND************************

.subckt AND N001 0 N003 N004 OUT
M1 N001 N003 N002 N001 pfet l=0.2u w=2u
M2 N001 N004 N002 N001 pfet l=0.2u w=2u
M3 N002 N003 N005 0 nfet l=0.2u w=1u
M5 N001 N002 OUT N001 pfet l=0.2u w=2u
M6 OUT N002 0 0 nfet l=0.2u w=1u
M4 N005 N004 0 0 nfet l=0.2u w=1u
.ends AND


****************OR************************

.subckt OR 1_d 0 v_a v_b OR
M1 1_d v_a N003 1_d pfet l=0.2u w=0.24u
M2 N003 v_b N005 1_d pfet l=0.2u w=0.24u
M3 1_d N005 OR 1_d pfet l=0.2u w=0.24u
M4 N005 v_a 0 0 nfet l=0.2u w=0.24u
M5 N005 v_b 0 0 nfet l=0.2u w=0.24u
M6 OR N005 0 0 nfet l=0.2u w=0.24u
.ends OR


****************clkDivider_50%_*********************

XU1 0 1_d N004 0 0 Q0 N004 clk DFFSR
XU2 0 1_d N005 0 0 Q1 N005 N004 DFFSR
XU3 0 1_d N006 0 0 Q2 N006 N005 DFFSR
XU4 0 1_d N007 0 N003 Q3 N007 Q2 DFFSR
XU5 0 1_d N008 0 N003 clk1 N008 N007 DFFSR
XU6 1_d 0 Q3 clk1 N003 AND
XU7 0 1_d clk1 0 0 N002 NC_11 N006 DFFSR
XU8 1_d 0 clk1 N002 clk_out OR


****************************************************

V1 clk 0 PULSE(0 1.8 1n 1n 1n 0.25u 0.5u)
V2 1_d 0 1.8

****************************************************

.tran 20us

*.lib C:\Users\ananya\Desktop\OR.cir
*.lib C:\Users\ananya\Documents\LTspiceXVII\active_high_with_qbar.cir
*.lib E:\VSD_Internship\progress\CIR files\ANDnew.cir

*.control
*run
*plot V(clk_out) V(clk)
*.endc
.end
